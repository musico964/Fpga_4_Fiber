-- megafunction wizard: %ALTGX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: alt2gxb 

-- ============================================================
-- File Name: gxb_transceiver.vhd
-- Megafunction Name(s):
-- 			alt2gxb
--
-- Simulation Library Files(s):
-- 			stratixiigx_hssi;sgate
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


-- related_files : gxb_transceiver.vhd
-- ipfs_files : gxb_transceiver.vho

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY gxb_transceiver IS
	PORT
	(
		cal_blk_clk		: IN STD_LOGIC ;
		pll_inclk		: IN STD_LOGIC ;
		rx_analogreset		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		rx_datain		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		rx_digitalreset		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		rx_enapatternalign		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		tx_ctrlenable		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		tx_datain		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		tx_digitalreset		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		pll_locked		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		rx_clkout		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		rx_ctrldetect		: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		rx_dataout		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		rx_disperr		: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		rx_errdetect		: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		rx_freqlocked		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		rx_patterndetect		: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		rx_syncstatus		: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		tx_clkout		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		tx_dataout		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0)
	);
END gxb_transceiver;


ARCHITECTURE SYN OF gxb_transceiver IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire11_bv	: BIT_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (0 DOWNTO 0);



	COMPONENT alt2gxb
	GENERIC (
		cmu_pll_inclock_period		: NATURAL;
		cmu_pll_loop_filter_resistor_control		: NATURAL;
		digitalreset_port_width		: NATURAL;
		enable_pll_inclk_alt_drive_rx_cru		: STRING;
		enable_pll_inclk_drive_rx_cru		: STRING;
		en_local_clk_div_ctrl		: STRING;
		equalizer_ctrl_a_setting		: NATURAL;
		equalizer_ctrl_b_setting		: NATURAL;
		equalizer_ctrl_c_setting		: NATURAL;
		equalizer_ctrl_d_setting		: NATURAL;
		equalizer_ctrl_v_setting		: NATURAL;
		equalizer_dcgain_setting		: NATURAL;
		intended_device_family		: STRING;
		loopback_mode		: STRING;
		lpm_hint		: STRING;
		lpm_type		: STRING;
		number_of_channels		: NATURAL;
		operation_mode		: STRING;
		pll_legal_multiplier_list		: STRING;
		preemphasis_ctrl_1stposttap_setting		: NATURAL;
		preemphasis_ctrl_2ndposttap_inv_setting		: STRING;
		preemphasis_ctrl_2ndposttap_setting		: NATURAL;
		preemphasis_ctrl_pretap_inv_setting		: STRING;
		preemphasis_ctrl_pretap_setting		: NATURAL;
		protocol		: STRING;
		receiver_termination		: STRING;
		reconfig_dprio_mode		: NATURAL;
		reverse_loopback_mode		: STRING;
		rx_8b_10b_compatibility_mode		: STRING;
		rx_8b_10b_mode		: STRING;
		rx_align_pattern		: STRING;
		rx_align_pattern_length		: NATURAL;
		rx_allow_align_polarity_inversion		: STRING;
		rx_allow_pipe_polarity_inversion		: STRING;
		rx_bandwidth_mode		: NATURAL;
		rx_bitslip_enable		: STRING;
		rx_byte_ordering_mode		: STRING;
		rx_channel_width		: NATURAL;
		rx_common_mode		: STRING;
		rx_cru_pre_divide_by		: NATURAL;
		rx_datapath_protocol		: STRING;
		rx_data_rate		: NATURAL;
		rx_data_rate_remainder		: NATURAL;
		rx_disable_auto_idle_insertion		: STRING;
		rx_enable_bit_reversal		: STRING;
		rx_enable_deep_align_byte_swap		: STRING;
		rx_enable_lock_to_data_sig		: STRING;
		rx_enable_lock_to_refclk_sig		: STRING;
		rx_enable_self_test_mode		: STRING;
		rx_enable_true_complement_match_in_word_align		: STRING;
		rx_flip_rx_out		: STRING;
		rx_force_signal_detect		: STRING;
		rx_ppmselect		: NATURAL;
		rx_rate_match_fifo_mode		: STRING;
		rx_run_length_enable		: STRING;
		rx_signal_detect_threshold		: NATURAL;
		rx_use_align_state_machine		: STRING;
		rx_use_clkout		: STRING;
		rx_use_coreclk		: STRING;
		rx_use_deserializer_double_data_mode		: STRING;
		rx_use_deskew_fifo		: STRING;
		rx_use_double_data_mode		: STRING;
		rx_use_rising_edge_triggered_pattern_align		: STRING;
		transmitter_termination		: STRING;
		tx_8b_10b_compatibility_mode		: STRING;
		tx_8b_10b_mode		: STRING;
		tx_allow_polarity_inversion		: STRING;
		tx_analog_power		: STRING;
		tx_channel_width		: NATURAL;
		tx_common_mode		: STRING;
		tx_data_rate		: NATURAL;
		tx_data_rate_remainder		: NATURAL;
		tx_enable_bit_reversal		: STRING;
		tx_enable_idle_selection		: STRING;
		tx_enable_self_test_mode		: STRING;
		tx_flip_tx_in		: STRING;
		tx_force_disparity_mode		: STRING;
		tx_refclk_divide_by		: NATURAL;
		tx_transmit_protocol		: STRING;
		tx_use_coreclk		: STRING;
		tx_use_double_data_mode		: STRING;
		tx_use_serializer_double_data_mode		: STRING;
		use_calibration_block		: STRING;
		vod_ctrl_setting		: NATURAL
	);
	PORT (
			pll_inclk	: IN STD_LOGIC ;
			rx_patterndetect	: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
			cal_blk_clk	: IN STD_LOGIC ;
			pll_locked	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_freqlocked	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_revbitorderwa	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_analogreset	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_datain	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_digitalreset	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_disperr	: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
			rx_enapatternalign	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_syncstatus	: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
			rx_clkout	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_ctrldetect	: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
			rx_dataout	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			rx_errdetect	: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
			tx_ctrlenable	: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
			tx_datain	: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			tx_digitalreset	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			tx_clkout	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			tx_dataout	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	sub_wire11_bv(0 DOWNTO 0) <= "0";
	sub_wire11    <= To_stdlogicvector(sub_wire11_bv);
	rx_patterndetect    <= sub_wire0(1 DOWNTO 0);
	pll_locked    <= sub_wire1(0 DOWNTO 0);
	rx_freqlocked    <= sub_wire2(0 DOWNTO 0);
	rx_disperr    <= sub_wire3(1 DOWNTO 0);
	rx_syncstatus    <= sub_wire4(1 DOWNTO 0);
	rx_clkout    <= sub_wire5(0 DOWNTO 0);
	rx_ctrldetect    <= sub_wire6(1 DOWNTO 0);
	rx_dataout    <= sub_wire7(15 DOWNTO 0);
	rx_errdetect    <= sub_wire8(1 DOWNTO 0);
	tx_clkout    <= sub_wire9(0 DOWNTO 0);
	tx_dataout    <= sub_wire10(0 DOWNTO 0);

	alt2gxb_component : alt2gxb
	GENERIC MAP (
		cmu_pll_inclock_period => 16000,
		cmu_pll_loop_filter_resistor_control => 3,
		digitalreset_port_width => 1,
		enable_pll_inclk_alt_drive_rx_cru => "true",
		enable_pll_inclk_drive_rx_cru => "true",
		en_local_clk_div_ctrl => "true",
		equalizer_ctrl_a_setting => 0,
		equalizer_ctrl_b_setting => 0,
		equalizer_ctrl_c_setting => 0,
		equalizer_ctrl_d_setting => 0,
		equalizer_ctrl_v_setting => 0,
		equalizer_dcgain_setting => 0,
		intended_device_family => "Arria GX",
		loopback_mode => "none",
		lpm_hint => "CBX_MODULE_PREFIX=gxb_transceiver",
		lpm_type => "alt2gxb",
		number_of_channels => 1,
		operation_mode => "duplex",
		pll_legal_multiplier_list => "disable_4_5_mult_above_3125",
		preemphasis_ctrl_1stposttap_setting => 0,
		preemphasis_ctrl_2ndposttap_inv_setting => "false",
		preemphasis_ctrl_2ndposttap_setting => 0,
		preemphasis_ctrl_pretap_inv_setting => "false",
		preemphasis_ctrl_pretap_setting => 0,
		protocol => "3g_basic",
		receiver_termination => "oct_100_ohms",
		reconfig_dprio_mode => 0,
		reverse_loopback_mode => "none",
		rx_8b_10b_compatibility_mode => "true",
		rx_8b_10b_mode => "normal",
		rx_align_pattern => "0101111100",
		rx_align_pattern_length => 10,
		rx_allow_align_polarity_inversion => "false",
		rx_allow_pipe_polarity_inversion => "false",
		rx_bandwidth_mode => 1,
		rx_bitslip_enable => "false",
		rx_byte_ordering_mode => "none",
		rx_channel_width => 16,
		rx_common_mode => "0.9v",
		rx_cru_pre_divide_by => 1,
		rx_datapath_protocol => "basic",
		rx_data_rate => 2500,
		rx_data_rate_remainder => 0,
		rx_disable_auto_idle_insertion => "false",
		rx_enable_bit_reversal => "false",
		rx_enable_deep_align_byte_swap => "false",
		rx_enable_lock_to_data_sig => "false",
		rx_enable_lock_to_refclk_sig => "false",
		rx_enable_self_test_mode => "false",
		rx_enable_true_complement_match_in_word_align => "false",
		rx_flip_rx_out => "false",
		rx_force_signal_detect => "true",
		rx_ppmselect => 1,
		rx_rate_match_fifo_mode => "none",
		rx_run_length_enable => "false",
		rx_signal_detect_threshold => 2,
		rx_use_align_state_machine => "false",
		rx_use_clkout => "true",
		rx_use_coreclk => "false",
		rx_use_deserializer_double_data_mode => "false",
		rx_use_deskew_fifo => "false",
		rx_use_double_data_mode => "true",
		rx_use_rising_edge_triggered_pattern_align => "false",
		transmitter_termination => "oct_100_ohms",
		tx_8b_10b_compatibility_mode => "true",
		tx_8b_10b_mode => "normal",
		tx_allow_polarity_inversion => "false",
		tx_analog_power => "1.5v",
		tx_channel_width => 16,
		tx_common_mode => "0.6v",
		tx_data_rate => 2500,
		tx_data_rate_remainder => 0,
		tx_enable_bit_reversal => "false",
		tx_enable_idle_selection => "false",
		tx_enable_self_test_mode => "false",
		tx_flip_tx_in => "false",
		tx_force_disparity_mode => "false",
		tx_refclk_divide_by => 1,
		tx_transmit_protocol => "basic",
		tx_use_coreclk => "false",
		tx_use_double_data_mode => "true",
		tx_use_serializer_double_data_mode => "false",
		use_calibration_block => "true",
		vod_ctrl_setting => 3
	)
	PORT MAP (
		pll_inclk => pll_inclk,
		cal_blk_clk => cal_blk_clk,
		rx_revbitorderwa => sub_wire11,
		rx_analogreset => rx_analogreset,
		rx_datain => rx_datain,
		rx_digitalreset => rx_digitalreset,
		rx_enapatternalign => rx_enapatternalign,
		tx_ctrlenable => tx_ctrlenable,
		tx_datain => tx_datain,
		tx_digitalreset => tx_digitalreset,
		rx_patterndetect => sub_wire0,
		pll_locked => sub_wire1,
		rx_freqlocked => sub_wire2,
		rx_disperr => sub_wire3,
		rx_syncstatus => sub_wire4,
		rx_clkout => sub_wire5,
		rx_ctrldetect => sub_wire6,
		rx_dataout => sub_wire7,
		rx_errdetect => sub_wire8,
		tx_clkout => sub_wire9,
		tx_dataout => sub_wire10
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ALT_SIMLIB_GEN STRING "1"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria GX"
-- Retrieval info: PRIVATE: NUM_KEYS NUMERIC "30"
-- Retrieval info: PRIVATE: RECONFIG_PROTOCOL STRING "BASIC"
-- Retrieval info: PRIVATE: RECONFIG_SUBPROTOCOL STRING "none"
-- Retrieval info: PRIVATE: RX_ENABLE_DC_COUPLING STRING "false"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WIZ_DATA_RATE STRING "2500"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INCLK_FREQ_ARRAY STRING "100 100"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A STRING "2000"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A_UNIT STRING "Mbps"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B STRING "100"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B_UNIT STRING "MHz"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_SELECTION NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_FREQ STRING "62.5"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_ENABLE_EQUALIZER_CTRL NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_EQUALIZER_CTRL_SETTING NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_FORCE_DEFAULT_SETTINGS NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_INCLK_FREQ STRING "62.5"
-- Retrieval info: PRIVATE: WIZ_INCLK_FREQ_ARRAY STRING "50.0 62.5 78.125 100.0 125.0 156.25 250.0 312.5 500.0"
-- Retrieval info: PRIVATE: WIZ_INPUT_A STRING "2500"
-- Retrieval info: PRIVATE: WIZ_INPUT_A_UNIT STRING "Mbps"
-- Retrieval info: PRIVATE: WIZ_INPUT_B STRING "62.5"
-- Retrieval info: PRIVATE: WIZ_INPUT_B_UNIT STRING "MHz"
-- Retrieval info: PRIVATE: WIZ_INPUT_SELECTION NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_SUBPROTOCOL STRING "No Loopback"
-- Retrieval info: PRIVATE: WIZ_WORD_ALIGN_FLIP_PATTERN STRING "0"
-- Retrieval info: CONSTANT: CMU_PLL_INCLOCK_PERIOD NUMERIC "16000"
-- Retrieval info: CONSTANT: CMU_PLL_LOOP_FILTER_RESISTOR_CONTROL NUMERIC "3"
-- Retrieval info: CONSTANT: DIGITALRESET_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: ENABLE_PLL_INCLK_ALT_DRIVE_RX_CRU STRING "true"
-- Retrieval info: CONSTANT: ENABLE_PLL_INCLK_DRIVE_RX_CRU STRING "true"
-- Retrieval info: CONSTANT: EN_LOCAL_CLK_DIV_CTRL STRING "true"
-- Retrieval info: CONSTANT: EQUALIZER_CTRL_A_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: EQUALIZER_CTRL_B_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: EQUALIZER_CTRL_C_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: EQUALIZER_CTRL_D_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: EQUALIZER_CTRL_V_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: EQUALIZER_DCGAIN_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Arria GX"
-- Retrieval info: CONSTANT: LOOPBACK_MODE STRING "none"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "alt2gxb"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "1"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "duplex"
-- Retrieval info: CONSTANT: PLL_LEGAL_MULTIPLIER_LIST STRING "disable_4_5_mult_above_3125"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_1STPOSTTAP_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_2NDPOSTTAP_INV_SETTING STRING "false"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_2NDPOSTTAP_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_PRETAP_INV_SETTING STRING "false"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_PRETAP_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: PROTOCOL STRING "3g_basic"
-- Retrieval info: CONSTANT: RECEIVER_TERMINATION STRING "oct_100_ohms"
-- Retrieval info: CONSTANT: RECONFIG_DPRIO_MODE NUMERIC "0"
-- Retrieval info: CONSTANT: REVERSE_LOOPBACK_MODE STRING "none"
-- Retrieval info: CONSTANT: RX_8B_10B_COMPATIBILITY_MODE STRING "true"
-- Retrieval info: CONSTANT: RX_8B_10B_MODE STRING "normal"
-- Retrieval info: CONSTANT: RX_ALIGN_PATTERN STRING "0101111100"
-- Retrieval info: CONSTANT: RX_ALIGN_PATTERN_LENGTH NUMERIC "10"
-- Retrieval info: CONSTANT: RX_ALLOW_ALIGN_POLARITY_INVERSION STRING "false"
-- Retrieval info: CONSTANT: RX_ALLOW_PIPE_POLARITY_INVERSION STRING "false"
-- Retrieval info: CONSTANT: RX_BANDWIDTH_MODE NUMERIC "1"
-- Retrieval info: CONSTANT: RX_BITSLIP_ENABLE STRING "false"
-- Retrieval info: CONSTANT: RX_BYTE_ORDERING_MODE STRING "none"
-- Retrieval info: CONSTANT: RX_CHANNEL_WIDTH NUMERIC "16"
-- Retrieval info: CONSTANT: RX_COMMON_MODE STRING "0.9v"
-- Retrieval info: CONSTANT: RX_CRU_PRE_DIVIDE_BY NUMERIC "1"
-- Retrieval info: CONSTANT: RX_DATAPATH_PROTOCOL STRING "basic"
-- Retrieval info: CONSTANT: RX_DATA_RATE NUMERIC "2500"
-- Retrieval info: CONSTANT: RX_DATA_RATE_REMAINDER NUMERIC "0"
-- Retrieval info: CONSTANT: RX_DISABLE_AUTO_IDLE_INSERTION STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_BIT_REVERSAL STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_DEEP_ALIGN_BYTE_SWAP STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_LOCK_TO_DATA_SIG STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_LOCK_TO_REFCLK_SIG STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_SELF_TEST_MODE STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_TRUE_COMPLEMENT_MATCH_IN_WORD_ALIGN STRING "false"
-- Retrieval info: CONSTANT: RX_FLIP_RX_OUT STRING "false"
-- Retrieval info: CONSTANT: RX_FORCE_SIGNAL_DETECT STRING "true"
-- Retrieval info: CONSTANT: RX_PPMSELECT NUMERIC "1"
-- Retrieval info: CONSTANT: RX_RATE_MATCH_FIFO_MODE STRING "none"
-- Retrieval info: CONSTANT: RX_RUN_LENGTH_ENABLE STRING "false"
-- Retrieval info: CONSTANT: RX_SIGNAL_DETECT_THRESHOLD NUMERIC "2"
-- Retrieval info: CONSTANT: RX_USE_ALIGN_STATE_MACHINE STRING "false"
-- Retrieval info: CONSTANT: RX_USE_CLKOUT STRING "true"
-- Retrieval info: CONSTANT: RX_USE_CORECLK STRING "false"
-- Retrieval info: CONSTANT: RX_USE_DESERIALIZER_DOUBLE_DATA_MODE STRING "false"
-- Retrieval info: CONSTANT: RX_USE_DESKEW_FIFO STRING "false"
-- Retrieval info: CONSTANT: RX_USE_DOUBLE_DATA_MODE STRING "true"
-- Retrieval info: CONSTANT: RX_USE_RISING_EDGE_TRIGGERED_PATTERN_ALIGN STRING "false"
-- Retrieval info: CONSTANT: TRANSMITTER_TERMINATION STRING "oct_100_ohms"
-- Retrieval info: CONSTANT: TX_8B_10B_COMPATIBILITY_MODE STRING "true"
-- Retrieval info: CONSTANT: TX_8B_10B_MODE STRING "normal"
-- Retrieval info: CONSTANT: TX_ALLOW_POLARITY_INVERSION STRING "false"
-- Retrieval info: CONSTANT: TX_ANALOG_POWER STRING "1.5v"
-- Retrieval info: CONSTANT: TX_CHANNEL_WIDTH NUMERIC "16"
-- Retrieval info: CONSTANT: TX_COMMON_MODE STRING "0.6v"
-- Retrieval info: CONSTANT: TX_DATA_RATE NUMERIC "2500"
-- Retrieval info: CONSTANT: TX_DATA_RATE_REMAINDER NUMERIC "0"
-- Retrieval info: CONSTANT: TX_ENABLE_BIT_REVERSAL STRING "false"
-- Retrieval info: CONSTANT: TX_ENABLE_IDLE_SELECTION STRING "false"
-- Retrieval info: CONSTANT: TX_ENABLE_SELF_TEST_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_FLIP_TX_IN STRING "false"
-- Retrieval info: CONSTANT: TX_FORCE_DISPARITY_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_REFCLK_DIVIDE_BY NUMERIC "1"
-- Retrieval info: CONSTANT: TX_TRANSMIT_PROTOCOL STRING "basic"
-- Retrieval info: CONSTANT: TX_USE_CORECLK STRING "false"
-- Retrieval info: CONSTANT: TX_USE_DOUBLE_DATA_MODE STRING "true"
-- Retrieval info: CONSTANT: TX_USE_SERIALIZER_DOUBLE_DATA_MODE STRING "false"
-- Retrieval info: CONSTANT: USE_CALIBRATION_BLOCK STRING "true"
-- Retrieval info: CONSTANT: VOD_CTRL_SETTING NUMERIC "3"
-- Retrieval info: USED_PORT: cal_blk_clk 0 0 0 0 INPUT NODEFVAL "cal_blk_clk"
-- Retrieval info: USED_PORT: pll_inclk 0 0 0 0 INPUT NODEFVAL "pll_inclk"
-- Retrieval info: USED_PORT: pll_locked 0 0 1 0 OUTPUT NODEFVAL "pll_locked[0..0]"
-- Retrieval info: USED_PORT: rx_analogreset 0 0 1 0 INPUT NODEFVAL "rx_analogreset[0..0]"
-- Retrieval info: USED_PORT: rx_clkout 0 0 1 0 OUTPUT NODEFVAL "rx_clkout[0..0]"
-- Retrieval info: USED_PORT: rx_ctrldetect 0 0 2 0 OUTPUT NODEFVAL "rx_ctrldetect[1..0]"
-- Retrieval info: USED_PORT: rx_datain 0 0 1 0 INPUT NODEFVAL "rx_datain[0..0]"
-- Retrieval info: USED_PORT: rx_dataout 0 0 16 0 OUTPUT NODEFVAL "rx_dataout[15..0]"
-- Retrieval info: USED_PORT: rx_digitalreset 0 0 1 0 INPUT NODEFVAL "rx_digitalreset[0..0]"
-- Retrieval info: USED_PORT: rx_disperr 0 0 2 0 OUTPUT NODEFVAL "rx_disperr[1..0]"
-- Retrieval info: USED_PORT: rx_enapatternalign 0 0 1 0 INPUT NODEFVAL "rx_enapatternalign[0..0]"
-- Retrieval info: USED_PORT: rx_errdetect 0 0 2 0 OUTPUT NODEFVAL "rx_errdetect[1..0]"
-- Retrieval info: USED_PORT: rx_freqlocked 0 0 1 0 OUTPUT NODEFVAL "rx_freqlocked[0..0]"
-- Retrieval info: USED_PORT: rx_patterndetect 0 0 2 0 OUTPUT NODEFVAL "rx_patterndetect[1..0]"
-- Retrieval info: USED_PORT: rx_syncstatus 0 0 2 0 OUTPUT NODEFVAL "rx_syncstatus[1..0]"
-- Retrieval info: USED_PORT: tx_clkout 0 0 1 0 OUTPUT NODEFVAL "tx_clkout[0..0]"
-- Retrieval info: USED_PORT: tx_ctrlenable 0 0 2 0 INPUT NODEFVAL "tx_ctrlenable[1..0]"
-- Retrieval info: USED_PORT: tx_datain 0 0 16 0 INPUT NODEFVAL "tx_datain[15..0]"
-- Retrieval info: USED_PORT: tx_dataout 0 0 1 0 OUTPUT NODEFVAL "tx_dataout[0..0]"
-- Retrieval info: USED_PORT: tx_digitalreset 0 0 1 0 INPUT NODEFVAL "tx_digitalreset[0..0]"
-- Retrieval info: CONNECT: @cal_blk_clk 0 0 0 0 cal_blk_clk 0 0 0 0
-- Retrieval info: CONNECT: @pll_inclk 0 0 0 0 pll_inclk 0 0 0 0
-- Retrieval info: CONNECT: @rx_analogreset 0 0 1 0 rx_analogreset 0 0 1 0
-- Retrieval info: CONNECT: @rx_datain 0 0 1 0 rx_datain 0 0 1 0
-- Retrieval info: CONNECT: @rx_digitalreset 0 0 1 0 rx_digitalreset 0 0 1 0
-- Retrieval info: CONNECT: @rx_enapatternalign 0 0 1 0 rx_enapatternalign 0 0 1 0
-- Retrieval info: CONNECT: @rx_revbitorderwa 0 0 1 0 GND 0 0 1 0
-- Retrieval info: CONNECT: @tx_ctrlenable 0 0 2 0 tx_ctrlenable 0 0 2 0
-- Retrieval info: CONNECT: @tx_datain 0 0 16 0 tx_datain 0 0 16 0
-- Retrieval info: CONNECT: @tx_digitalreset 0 0 1 0 tx_digitalreset 0 0 1 0
-- Retrieval info: CONNECT: pll_locked 0 0 1 0 @pll_locked 0 0 1 0
-- Retrieval info: CONNECT: rx_clkout 0 0 1 0 @rx_clkout 0 0 1 0
-- Retrieval info: CONNECT: rx_ctrldetect 0 0 2 0 @rx_ctrldetect 0 0 2 0
-- Retrieval info: CONNECT: rx_dataout 0 0 16 0 @rx_dataout 0 0 16 0
-- Retrieval info: CONNECT: rx_disperr 0 0 2 0 @rx_disperr 0 0 2 0
-- Retrieval info: CONNECT: rx_errdetect 0 0 2 0 @rx_errdetect 0 0 2 0
-- Retrieval info: CONNECT: rx_freqlocked 0 0 1 0 @rx_freqlocked 0 0 1 0
-- Retrieval info: CONNECT: rx_patterndetect 0 0 2 0 @rx_patterndetect 0 0 2 0
-- Retrieval info: CONNECT: rx_syncstatus 0 0 2 0 @rx_syncstatus 0 0 2 0
-- Retrieval info: CONNECT: tx_clkout 0 0 1 0 @tx_clkout 0 0 1 0
-- Retrieval info: CONNECT: tx_dataout 0 0 1 0 @tx_dataout 0 0 1 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL gxb_transceiver.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL gxb_transceiver.ppf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL gxb_transceiver.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL gxb_transceiver.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL gxb_transceiver.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL gxb_transceiver_inst.vhd FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL gxb_transceiver.vho TRUE
-- Retrieval info: LIB_FILE: stratixiigx_hssi
-- Retrieval info: LIB_FILE: sgate
-- Retrieval info: CBX_MODULE_PREFIX: ON
